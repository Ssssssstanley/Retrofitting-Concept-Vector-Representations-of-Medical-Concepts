CUI1	CUI2	Mean
C0017601	C0232197	279
C0006949	C0031507	370.5
C0878544	C0000970	241
C0019340	C0020550	142.5
C0036494	C0027497	870.75
C0009186	C0019655	981.25
C0002962	C0070166	673.75
C0061851	C0022046	294.25
C0036572	C0021641	332.75
C0036690	C0013404	434.5
C0028738	C0021167	365.75
C0036494	C0001962	465
C0013456	C0034880	760.25
C0032064	C0008402	255.25
C0001367	C0209227	1052
C0027497	C0027498	1039.25
C0162275	C0159075	334.5
C0009951	C0001962	835.25
C0242723	C0024530	1239.25
C0033687	C0011847	1047
C0017160	C0086073	391
C0020639	C0020175	519.75
C0213771	C0073992	1118.5
C0162275	C0016410	383
C0021641	C0017687	448.75
C0086543	C0043144	217.25
C0025605	C0040610	663.5
C0011847	C0033860	412
C0948786	C0030232	1180.75
C0232471	C0016860	935.25
C0031763	C0003564	284.25
C0032617	C0159075	189.5
C0033860	C0025287	222.25
C0042755	C0013132	543
C0009421	C0019158	565
C0917801	C0085631	882.5
C0442874	C0025598	487.75
C0033860	C0003864	1148.75
C0041296	C0149651	631.25
C0028754	C0011847	1142.25
C0040038	C0019079	852
C0032285	C0007561	867.25
C0114873	C0076107	716.25
C0086543	C0025598	272.75
C1623038	C0301532	523
C0036572	C0006949	798
C0086543	C0021641	391
C0002871	C0206160	897
C0009951	C0006949	844
C0029456	C0032950	755
C0036572	C0031507	1001.75
C0885057	C0016157	933.75
C0242339	C0016157	921.5
C0232197	C0002962	725.5
C0007557	C0007561	1154.5
C0011053	C0004134	582.75
C0220892	C0007546	1078.75
C0011847	C0021641	1155.25
C0018995	C0003126	382
C0022116	C0152149	398
C0030232	C0004057	406.75
C0013456	C0233212	367.75
C0019340	C0008370	475.25
C0242339	C0008402	889.5
C0034494	C0702166	256.25
C0032064	C0001416	816.25
C0159075	C0232955	239
C0001975	C0012772	743
C0009214	C0027358	578.5
C0043031	C0004057	1019.75
C0042313	C0017642	829.25
C0009187	C0025289	791.25
C0030232	C0043031	638.25
C0002940	C0029456	231.25
C0022116	C0025859	823.75
C0016204	C0017687	727.5
C0007546	C0007716	1323
C0029456	C0087086	240.75
C0014038	C0025289	1037.75
C0684275	C0040038	450
C0003864	C0003862	1091
C0152447	C0040822	342.5
C0003128	C0079083	662.75
C0001924	C0019134	377.5
C0032617	C0021641	766.75
C0037384	C0038450	492.75
C0033860	C0054836	194.75
C0019112	C0021359	191.25
C0014544	C0031412	940.75
C0014544	C0001975	566.75
C0033860	C0037763	221.25
C0037384	C0023992	242
C0003850	C0008402	510.25
C0854467	C0037384	358
C0032285	C0036690	959.25
C0019270	C0497327	237.75
C0018926	C0027498	1012.25
C0003862	C0030193	1206.25
C0040165	C0023660	270.25
C0032285	C0013404	833.75
C0741439	C0025287	776.75
C0017601	C0232197	276
C0036494	C0007297	893.25
C0003862	C0149651	317.5
C0684275	C0017642	169
C0013428	C0070166	212.5
C0231236	C0042755	294.5
C0002940	C0947651	340.5
C0009262	C0032950	851.25
C0019270	C0006982	418
C1257763	C0036572	396.5
C0086543	C0030305	307.5
C0001962	C0001975	1265.5
C0020550	C0036572	792.25
C0116569	C0002598	1058.75
C0021359	C0079083	853.5
C0003862	C0027796	763.5
C0003129	C0033487	477.75
C0012833	C0004147	617.75
C0030305	C0021641	749.5
C0017160	C0021641	351.75
C0023530	C0007537	343
C0019655	C0032950	290
C0442874	C0009806	477.25
C0149651	C0013404	930.75
C0018991	C0070166	704.5
C0026946	C0286651	300.5
C0035435	C0009262	775.25
C0013404	C0220892	384
C1623038	C0018926	1040.25
C0877781	C0018681	748.75
C0023992	C0005632	767
C0920289	C0015672	1186.5
C0878544	C0039070	869.5
C0003129	C0036572	748
C0036494	C0001962	646
C0242339	C0060277	239
C0039730	C0040822	231.5
C0009951	C0085208	869.25
C0002962	C0028351	398.75
C0027121	C0025815	792.75
C0003128	C0152149	558.25
C0013456	C0002645	855.25
C0022116	C0995182	253.5
C0006277	C0298130	737.25
C0286651	C0024027	1174.75
C0032285	C1883552	633.75
C0037763	C0016860	415.75
C0040485	C0014806	343
C0011603	C1998461	1188
C0947651	C0022614	293.75
C0003850	C0022116	751.75
C0018995	C0032617	309.5
C0025587	C0040460	573.25
C0011175	C0038187	977
C0009319	C0014544	163
C0011847	C0085602	1031.5
C0162275	C0038187	1225.25
C0036572	C0042291	911
C0018081	C0070166	173
C0301532	C0039840	893
C0020676	C1883552	904.75
C0039730	C0019045	1307
C0206160	C0004057	670.75
C0026946	C0079083	340.5
C0026946	C0025289	975.5
C0030232	C0060277	901.75
C0332566	C0332573	1090
C0018834	C0020740	644
C0995182	C0020264	187.5
C0009214	C0011816	830.75
C0001047	C0001443	256.25
C0086073	C0032950	856
C0037763	C0151818	665.75
C0011991	C0007537	508.75
C0007559	C0007561	1086.5
C0030193	C0026549	996.75
C0027358	C0015846	484.25
C0042384	C0018991	363.5
C0009262	C0033209	1098.75
C0126174	C0216784	1243.5
C1623038	C0002871	727.5
C0055003	C0004899	648.25
C0037354	C0042214	721.5
C0038187	C0152149	145.5
C0031763	C0011603	957.75
C0011777	C0246719	472
C0019158	C0000970	880.25
C0022116	C0013132	468.75
C0019270	C0013456	179.75
C0018021	C0011644	394
C0004134	C0001962	840.25
C0043528	C0004576	1136.75
C0035508	C0034642	1075.5
C0557875	C0004147	537
C0004153	C0002962	936
C0019158	C0018926	778
C0027358	C0026549	571.5
C0011991	C0009262	794.5
C0027121	C0026848	1103
C0006277	C0023992	242.75
C0013428	C0008809	615.5
C0282386	C0536495	1120.25
C0034880	C0005740	607.5
C0008168	C0007561	652.75
C0007537	C0007557	1174.5
C0014806	C0023660	430
C0020676	C0021359	598
C0081876	C0006681	971.75
C0007398	C0023380	890
C0036323	C0114873	201.75
C0085602	C0032617	1135.5
C1623038	C0286651	390.5
C0038450	C0037384	646.5
C0004147	C0016860	708.25
C0242453	C0008809	744.5
C0011175	C0013369	925.75
C0014025	C0065374	1280
C0235250	C0079083	765.25
C0206160	C0018926	427
C0041948	C0751229	657.5
C0026848	C0234369	555.25
C0021359	C0232197	346
C0162275	C0021641	891.5
C0005716	C0036572	579.75
C0006840	C0392071	383.5
C0019134	C0033603	691
C0878544	C0034642	705.75
C0026946	C0030193	355.25
C0033687	C0026196	285.25
C0002962	C0013404	642.25
C0004610	C0376288	445
C0242339	C0286651	1029.5
C0041948	C0013911	499.5
C0029456	C0878544	295.25
C0235250	C0027497	1240.25
C0242723	C0858529	331
C0442874	C0021641	754.75
C0036494	C0149651	306.25
C0060277	C0060277	1395
C0858529	C0023992	279.5
C0035435	C0000970	923.5
C0006309	C0043528	1195.75
C0004147	C0025859	1279.25
C0013911	C0006625	1290.25
C0003564	C0152149	214.25
C0038187	C0003123	1176.75
C0005747	C0043031	207.75
C0002680	C0002645	1238
C0002962	C0011991	270.75
C0016860	C0024730	658.5
C0041948	C0553735	551
C0021167	C0016860	739.5
C0040038	C0019134	969.75
C0015300	C0242453	243.5
C0041948	C0004057	256
C0006982	C0018242	240.25
C1998461	C0004899	203
C0019270	C0018021	354.75
C0011175	C0039070	897.75
C0231851	C0032617	303.25
C0003864	C0035435	1153.25
C0021359	C0003128	1192.75
C0006277	C0073992	939.25
C0026946	C0019655	1282.5
C0086543	C0011847	652.75
C1257763	C0162429	160.75
C0009951	C0014544	1302.75
C0010520	C0016410	365.5
C0021359	C0005747	225.25
C0442874	C0011847	1032
C0014806	C0002144	345.5
C0018834	C0081876	981.5
C0030232	C1883552	1109.5
C0231451	C0017245	258.75
C1883552	C0030552	1158.25
C0020676	C0040165	984.75
C0239779	C0221169	634
C0015300	C0040165	928.5
C0021359	C0003128	1276.5
C0012833	C0042571	1287
C0242339	C0002962	806
C0017536	C0376286	422
C0036572	C0995182	167.75
C0074393	C0016365	1138.75
C0031154	C0004134	281.75
C0246719	C0102118	1276.5
C0003862	C0159075	201
C0149651	C0009806	167.75
C0070166	C0286651	895.5
C0014563	C0028351	394.5
C0009806	C0011991	161
C0003864	C1623038	618.5
C0025289	C0041296	871.25
C0012833	C0001962	893.25
C0086543	C0027358	263.5
C0085631	C0026549	527.5
C0003126	C0003564	845
C0013132	C0006982	662.75
C1623038	C0025677	706.25
C0017601	C0018681	841.25
C0039070	C1883552	737
C2004489	C0018834	1106.5
C0032143	C0038418	762.75
C0052796	C0008809	965
C0007398	C0027358	458
C0003862	C0000970	869.25
C0005747	C0270327	321.25
C0085635	C0018681	632
C0025289	C0018681	1221.25
C0017628	C0289313	1128.25
C0004153	C0858529	997.75
C0003126	C0231617	274.5
C0235250	C0061851	738.5
C0002962	C0231618	666.25
C0398623	C0019079	469.75
C0028754	C0076275	1007.25
C0017642	C0020740	330.5
C0004153	C0021400	257.75
C0231655	C0018520	233.5
C0019209	C0019214	1164.75
C0003126	C0012265	293
C0025289	C0042313	960.25
C0751229	C0037384	764
C0392071	C0008809	981.25
C0016204	C0018520	802.25
C0016382	C0060277	511.5
C0152149	C0003564	199.25
C0018995	C0003864	858.25
C0149651	C0042878	360.5
C0152149	C0040460	567.75
C0232471	C0020175	935.75
C0036396	C0020740	854.5
C0006277	C0032285	1019.75
C0006840	C0025815	390.25
C0037384	C0001962	706.25
C0232197	C0357929	256
C0012265	C0012373	1045
C0002333	C0024002	1269
C0019158	C1623038	1173
C0013404	C0025815	836
C0149651	C0885057	194
C0035435	C0917801	384.75
C0035435	C0032950	883.25
C0011847	C0020456	1234.75
C0232197	C0043031	1106.75
C0877781	C0017887	298.75
C0040038	C0232197	1026.5
C0019079	C0043031	936.75
C0029456	C0246719	811.25
C0004134	C0009806	309.25
C0026946	C0009187	1137.25
C0036396	C0231236	375.25
C0009014	C0025859	921.25
C0003615	C0007546	889.5
C0007561	C0007557	1202.25
C0877781	C0000970	619.5
C0070166	C0043031	1183.5
C0017160	C0013369	1255.75
C0014544	C0019209	208.25
C0020639	C0020175	886.5
C0013404	C0073992	815.25
C0028978	C0025598	305.75
C0008838	C0061851	645.5
C0025815	C0032950	1387.5
C0022116	C0286651	953.25
C0231655	C0017887	246.75
C0026946	C0005716	1118.5
C0027497	C0061851	974
C0008402	C1142985	1184
C1883552	C0074554	889.75
C0152447	C0003564	233.25
C0079083	C0008838	1273.5
C0442874	C0039128	1034
C0039128	C0220892	1094.25
C0022251	C0025859	1031.5
C0027697	C0553735	807.5
C0013090	C0220892	680.75
C0041948	C0020740	393.25
C0034642	C0010520	687.5
C0231451	C0020175	338
C0152149	C0246719	307.5
C1623038	C0018995	956
C0030305	C0086543	342
C0030305	C0332566	348.5
C0040038	C0013404	962.5
C0019158	C0019209	910.25
C0034880	C0003564	431.75
C0040034	C0018834	328.5
C0003615	C0031154	934.75
C0025587	C0009262	792.25
C0741439	C1282609	683.25
C0028351	C0033487	784
C0035435	C0162323	1124.75
C0085593	C0037384	322.5
C0276185	C0752270	450
C1257763	C0010592	232.75
C0023530	C0005740	890
C0040165	C0279175	483.75
C0004153	C0152447	212.25
C0232197	C0040165	881.5
C0398623	C0043031	846.75
C0018991	C0018681	561.5
C0004153	C0040460	224.5
C0009024	C0037763	967
C0553735	C0027697	777.5
C0013404	C0027358	578.25
C0006309	C0027358	199.75
C0025287	C0020453	536.75
C0039730	C0060277	892.5
C0017887	C0025859	785.25
C1998461	C0025287	319.5
C0242706	C0076275	343.5
C0001882	C0029456	206.5
C0009806	C0012373	178.75
C0006840	C0026946	1151.25
C0074554	C0016157	923.5
C0009421	C0003129	668
C0002962	C0858529	863
C0042384	C0009951	372.5
C0039070	C0002333	618.25
C0018081	C0076275	193.75
C0242706	C0076275	197.25
C0036323	C0242723	1187.5
C0286651	C0074554	1330.75
C0037384	C0221232	327.5
C0003129	C0004134	496.75
C0009421	C0086543	265.25
C0085208	C0002600	309
C0003126	C0009806	244.25
C0018681	C0016382	413.25
C0741439	C0027497	503.25
C0031412	C0042291	1046.5
C0005740	C0012772	337.75
C0376286	C0038187	984.75
C0026946	C0025815	388.75
C0162323	C0003862	1126
C0878544	C0002962	861.5
C1623038	C0074554	498
C0020175	C0038187	1134.5
C0020676	C0009421	710.75
C0021400	C0002403	919
C0000970	C0020740	1067
C0242706	C0003129	252
C0022116	C0022251	837.5
C0003128	C0040485	228
C0041296	C0019079	789.5
C0232197	C0002962	788.5
C0020676	C0557875	948.75
C0039128	C0497327	960.5
C0079083	C0061851	940
C0013132	C0085593	395
C0003864	C0231236	333.25
C0011847	C0032617	1066
C0019079	C0018926	908.25
C0033687	C0065374	926.5
C0013132	C0023570	800.75
C0030232	C0001924	528.75
C0039128	C0018081	1132.25
C0086543	C0231655	288.5
C0014544	C0024002	836.5
C0001416	C0038450	666.25
C0018834	C0015620	893.5
C0149651	C0213771	846.75
C0004096	C0451641	286
C0040038	C0043031	964.75
C0232197	C0018520	348
C0178664	C0033687	858
C0028734	C0011847	775.25
C0036572	C0357929	190.75
C0231655	C0025587	870.25
C0002144	C0009262	1142.25
C0018995	C0003862	774.25
C0002403	C0874161	1193
C0025289	C0007561	1030
C0027121	C0286651	853.75
C0032285	C0010520	623.25
C0040038	C0039070	728.5
C0009090	C0017887	219.5
C0040034	C0003864	306.5
C0039070	C0004147	639.5
C0040822	C0023570	840.5
C0014544	C0003126	404.25
C0085631	C0040165	637.5
C0003128	C0013911	574
C0041834	C0031507	468.5
C0011175	C0006840	547
C0034642	C0034880	251.25
C0010137	C0001443	214.75
C0018681	C0000970	879.5
C0003864	C0025587	769
C0041834	C0040822	316
C0028754	C0037384	860
C0013404	C0010520	1052.25
C0041948	C0027497	621.25
C0242453	C0392071	964.75
C0019045	C0030193	505.25
C0009421	C0020456	922.25
C1883552	C0013911	956.25
C0232471	C0020175	819
C0013404	C0213771	1075.5
C0242339	C0032143	531.75
C0023530	C0220892	416.25
C0025289	C0025287	864.5
C1883552	C0017687	368
C0009806	C0042523	193
C0232197	C0004147	817.25
C0018021	C0042384	324.75
C0028734	C0004899	353.75
C0020550	C0029456	493.75
C0242339	C0020473	809.5
C0030232	C0948786	955
C0393080	C0016365	193.25
C0019079	C0033603	544
C0024902	C0013456	807.5
C0034642	C0016860	742
C0002871	C0043031	623.75
C0023570	C0006982	1533.5
C0011603	C0995182	695
C0009187	C0025815	388.5
C0557875	C0751229	1055.25
C0032617	C0162275	993.25
C0040460	C0004134	255.5
C0024730	C0000970	223
C0029877	C0025287	567
C0009024	C0085208	317.5
C0002871	C0070166	539.5
C0016157	C0074554	809.5
C0028734	C0001962	680.25
C1883552	C0010137	682
C0242339	C0009806	318.5
C0026946	C0242453	271.5
C0497327	C0995182	223.5
C0013369	C0116569	229.5
C0032064	C0006644	278.5
C0034494	C0947651	239
C0021400	C0032285	898.5
C0034494	C0234990	417.25
C0070166	C0021641	286.25
C0017536	C0233576	152.75
C0033860	C0004153	169.5
C0033497	C0085259	318.75
C0040460	C0076107	224.75
C0011633	C0026848	1019.5
C0038187	C0008838	319
C0003128	C0002453	1099.5
C0001824	C0002871	933.25
C0040485	C0037763	1104
C0557875	C0042523	233.75
C0357929	C0005740	227
C0018995	C0025023	212.25
C0003128	C0006982	326.25
C0231451	C0004899	261.25
C0001927	C0073992	949.5
C0003864	C0002726	724.25
C0010520	C0014563	456.5
C0015620	C0034665	1247.25
C0014544	C0022116	506.75
C0007297	C0027497	1168.75
C0232197	C0878544	764.5
C0043528	C0032064	997.25
C0025287	C0001367	713.5
C0000786	C0023860	781.5
C0013404	C0085631	593.25
C0014038	C0018681	1052.5
C0014544	C0246719	329.25
