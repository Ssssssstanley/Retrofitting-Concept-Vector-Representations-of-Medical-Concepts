CUI1	CUI2	Mean
C0878544	C0039070	794.75
C0086543	C0043144	499.25
C0018834	C0043066	1151.75
C0001927	C0298130	1165.5
C0041296	C0030232	869.5
C0231451	C0017245	732.75
C0231851	C0032617	527.25
C0031154	C0239779	804
C0040038	C0019079	778.25
C0003862	C0149651	917.5
C0007398	C0027358	753.5
C0043167	C0023343	827.75
C0003128	C0013911	535.25
C0442874	C0021641	1126.75
C1998461	C0004899	829.5
C0376286	C0038187	770.75
C0041834	C0040822	528
C0178664	C0033687	1061
C0032064	C0001416	753
C0001047	C0001443	586.5
C0004147	C0016860	895.5
C0011847	C0009214	615.75
C0086543	C0011847	1043
C0014806	C0002144	666.75
C1257763	C0162429	1070.25
C0041296	C0149651	865.75
C0019270	C0497327	570.25
C0020639	C0020175	957.25
C0019079	C0033603	798
C0042755	C0013132	663.75
C1623038	C0018926	1040
C0497327	C0033860	582.25
C0029456	C0087086	630.5
C0009806	C0011991	1023.5
C0116569	C0002598	695.75
C0002962	C0011991	553.5
C0000786	C0023860	1005.25
C0013404	C0027358	1064.5
C0013404	C0213771	1146.75
C0041948	C0553735	856.25
C0149651	C0013404	1070
C0039730	C0040822	678.5
C0037384	C0023992	699.75
C0030232	C0001924	987.5
C0020459	C0011847	1152
C0004153	C0022116	1170.5
C0004153	C0018834	618.5
C0029456	C0246719	771
C0011991	C0009262	947.25
C0013428	C0008809	1061
C0009421	C0003129	1099.5
C0013456	C1510450	1111.5
C0038450	C0037384	676.25
C0017887	C0025859	972.75
C0028738	C0021167	616.25
C0014544	C0006949	761
C0022251	C0025859	1064.25
C0017160	C0021641	668.25
C0018995	C0003862	899.25
C0029877	C0025287	848
C1623038	C0286651	1142.75
C0028734	C0001962	679.5
C0002962	C0018834	1139
C0013428	C0019079	593.5
C0001047	C0000970	1109
C0004093	C0006625	815.5
C0009024	C0037763	917
C0018995	C0003864	857.25
C0016204	C0018520	873
C0027358	C0026549	1189.25
C0239779	C0221169	1044.25
C0149651	C0009806	511.5
C0018991	C0070166	651.25
C0036396	C0231236	823.75
C0398623	C0043031	765.75
C0003128	C0152149	1006
C0020639	C0020175	710.5
C0021167	C0016860	779.75
C0014544	C0031412	1135.25
C0030305	C0011847	1063.75
C0014544	C0019209	747.75
C0017160	C0036572	785
C0149651	C0213771	1027
C1623038	C0019270	664
C0032617	C0021641	1085.5
C0011053	C0029877	1072.5
C0003864	C0231236	482.75
C0026848	C0234369	756
C0036494	C0001962	897
C0036572	C0085208	816.75
C0232197	C0040165	929.75
C0004134	C0009806	543.25
C0018021	C0011644	578.5
C0016293	C0012010	959.5
C0011175	C0006840	570.25
C0001416	C0038450	680.5
C0034642	C0010520	839
C0027358	C0015846	737
C0014544	C0001975	856.75
C0001367	C0209227	860.25
C0034880	C0005740	845.5
C0074554	C0016157	1119.75
C0041948	C0751229	806
C0398623	C0019079	717.75
C0332566	C0332573	943
C0162275	C0159075	704.75
C0040034	C0036396	443.5
C0030305	C0021641	1054.75
C0016410	C0014563	899.25
C0006840	C0025815	774.75
C0019079	C0043031	987.75
C0040485	C0014806	657.25
C0017160	C0086073	776
C0013404	C0220892	664
C0013404	C0025815	919.5
C0242723	C0858529	764.5
C0242723	C0025815	864.75
C0005716	C0036572	932
C0018681	C0016382	1002.25
C0032285	C0010520	1078.75
C0159075	C0232955	816.25
C0040038	C0011603	519.25
C0061851	C0022046	990
C0086543	C0021641	463.75
C0025815	C0032950	1180.25
C0025587	C0009262	742
C0009014	C0025859	884.5
C1883552	C0074554	726.25
C0009214	C0011816	1119.75
C0027121	C0026848	1049.75
C0032617	C0159075	964.75
C0022116	C0286651	971.25
C0002871	C0043031	926.5
C0246719	C0102118	850.25
C0086543	C0025598	573.75
C0885057	C0016157	824
C0009806	C0012373	508
C0021641	C0289313	990.25
C0242453	C0392071	1023
C0858529	C0023870	853.25
C0028754	C0076275	978.75
C0086073	C0032950	997.75
C0037384	C0038450	610
C0025605	C0040610	837.25
C0741439	C0027497	685.25
C0009951	C0085208	831
C0034880	C0003564	846.75
C0034494	C0234990	585
C0035435	C0009262	825.5
C0003128	C0040485	460.75
C0020676	C0009421	1033.75
C0004899	C0042313	1028.75
C0231451	C0020175	489.5
C0036572	C0006949	998.5
C0032064	C0006644	637
C0009187	C0025289	948
C0013911	C0079083	708.75
C0013090	C0220892	1109.5
C0014544	C0024002	469.25
C0014806	C0023660	688
C0086140	C0002658	597.5
C0041948	C0027497	974.5
C0013132	C0006982	943.5
C0553735	C0242453	867.5
C0025287	C0001367	989.5
C0043528	C0032064	1135
C0003128	C0006982	619.75
C0011847	C0032950	1099.5
C0013369	C0012833	1157
C0553735	C0027697	884.75
C0018995	C0032617	635.5
C0151818	C0036572	1058.5
C0948786	C0030232	1173.5
C0009421	C0086543	330.25
C0025587	C0040460	787.25
C0242706	C0003129	1059
C0231451	C0004899	474.25
C0025587	C0009014	774.75
C0040460	C0076107	518.75
C0042313	C0017642	824.75
C0005747	C0152149	588
C0024205	C0276185	612
C0026946	C0009187	1185.75
C0020550	C0036572	1121
C0004610	C0376288	698.5
C0085631	C0040165	943.75
C0014544	C0022116	477.5
C0282386	C0536495	1110.75
C0003615	C0007546	879.75
C0008168	C0007561	717.5
C0016382	C0060277	673.75
C0001924	C0019134	1011
C1623038	C0074554	1092.75
C0017536	C0376286	718.25
C0114873	C0076107	906
C1998461	C0025287	416.25
C0009187	C0025815	831.25
C0026946	C0030193	958.5
C0553735	C0013428	1064
C0085593	C0037384	650.75
C0011847	C0033860	787.5
C0085635	C0018681	1168.5
C0003126	C0231617	431.25
C0043066	C2004489	1179
C0231655	C0017887	732.25
C0231655	C0018520	505
C0006277	C0298130	702.5
C0035435	C0032950	720.5
C0026946	C0025815	550
C0017601	C0232197	528.5
C0392071	C0008809	1044.75
C0013132	C0085593	465
C0023530	C0005740	1036.5
C0023530	C0220892	640.25
C0035435	C0920289	833.5
C0206160	C0018926	487
C0271397	C1698636	1173
C0034494	C0947651	555.25
C0013428	C0152447	903.75
C0041834	C0031507	516.25
C0026946	C0286651	595.25
C0030232	C0004057	871.25
C0021641	C0017687	1261.5
C0038187	C0008838	788.25
C0026946	C0025289	812.25
C0007716	C0076275	564.25
C0301532	C0001975	1315.5
C0149651	C0042878	529.75
C0002940	C0947651	540.25
C0032285	C0025289	773
C0006309	C0043528	1214
C0011053	C0005747	438.75
C0702166	C0004134	343.5
C0009090	C0233576	669
C0031763	C0003564	441.25
C0019655	C0032950	789.5
C0014544	C0246719	818.5
C0086543	C0030305	473.5
C0398623	C0040038	1139
C0016157	C0074554	1276.5
C0001824	C0854467	1230.25
C0015300	C0019214	527.25
C0001975	C0012772	1244
C0004153	C0021400	416
C0006277	C0032285	1066.5
C0741439	C1282609	1174.5
C0040822	C0023570	1224.5
C0684275	C0017642	418.75
C0004905	C0012373	514.25
C0039730	C0019045	1218
C0019340	C0008370	525.75
C0002403	C0874161	1274.75
C0042523	C0752270	829.5
C0018081	C0076275	404.75
C0036494	C0007297	1233
C0011175	C0039070	1028.75
C0232471	C0020175	1249
C0009262	C0033209	1307.75
C0175848	C0043066	681.5
C0021359	C0005747	411.5
C0042384	C0018991	656.25
C0232471	C0016860	1171.75
C0020676	C1883552	1224.75
C0030552	C0221166	1253.25
C0032143	C0038418	899.5
C0010137	C0001443	409.75
C0877781	C0018681	1210.5
C0231236	C0042755	414.5
C0086543	C0014544	361
C0030232	C0948786	1248
C0034642	C0034880	409.5
C1257763	C0036572	488.5
C0878544	C0000970	417.25
C0013404	C0073992	843.5
C0917801	C0086140	475
C0242453	C0008809	815.5
C0019270	C0006982	462.5
C0020459	C0037384	444
C0013428	C0070166	415
C0006277	C0023992	582
C0041948	C0023870	582
C0036396	C0102118	446.5
C0036396	C0246719	473.5
C0006982	C0018242	746
C0036572	C0995182	392.5
C0003129	C0004134	444.75
C0017628	C0289313	1069.25
C0006277	C0073992	916
C0451641	C0002726	565.75
C0357929	C0005740	593.25
C0231655	C0025587	833.75
C0003126	C0009806	391
C0002962	C0014563	622.75
C0008350	C0006277	345
C0009024	C0085208	752
C0232197	C0087086	1285.75
C0009951	C0006949	1234.75
C0010592	C0032950	601.75
C0018021	C0020740	427.25
C0003862	C0717550	452.5
C0006840	C0026946	1161.25
C0010520	C0016410	420
C0858529	C0017887	1190
C0002871	C0206160	1187
C0026946	C0019655	1272.5
C0018546	C0004899	492.75
C0442874	C0039128	1225.75
C0242706	C0076275	564
C0557875	C0042523	603.75
C0276185	C0752270	531
C0033497	C0085259	500
C0017642	C0020740	601.25
C0033860	C0025287	470
C0009806	C0042523	662.5
C0019079	C0018926	1269.75
C0026946	C0242453	555.75
C0004134	C0022614	488.5
C0011603	C0995182	1286.25
C0242706	C0076275	446
C0042384	C0009951	438.75
C0011175	C0038187	1163.75
C0002333	C0024002	1034
C0878544	C0034642	1048.25
C0038187	C0152149	439.5
C0015300	C0242453	411.25
C0684275	C0019079	931.25
C0037763	C0036396	1068.25
C0004147	C0025859	1182.25
C0039730	C0060277	1199.25
C0242723	C0024530	1277
C0043528	C0004576	1270.25
C0023530	C0032285	722
C0003862	C0159075	670
C1998461	C0019134	1084.25
C0019270	C0018021	379.75
C0020676	C0009421	1197.25
C0004153	C0040460	455
C0741439	C0025287	1002.75
C0012833	C0015672	1231.25
C0152149	C0003564	448.5
C0947651	C0022614	752.5
C0021359	C0079083	1134.75
C0036396	C0020740	1054.25
C0162323	C0003862	1188.75
C0023413	C0025677	1111.25
C0002962	C0028351	474.5
C0276185	C0043066	460.75
C0242339	C0032143	615.75
C0040165	C0023660	365.25
C0040822	C0006982	1150.25
C0079083	C0008838	1303
C0152149	C0246719	448.25
C0995182	C0020264	399.75
C0041948	C0020740	482
C0003862	C0000970	1277
C0040165	C0279175	1071.25
C0017887	C0026549	1126
C0036572	C0357929	658.5
C0014544	C0003126	515.25
C1257763	C0010592	654.5
C0016860	C0024730	1093.5
C0086543	C0231655	460.75
C0003128	C0002453	1332
C0074393	C0016365	1350.5
C0016579	C0030554	641.75
C0018834	C0014724	560
C0001367	C0070122	604.75
C0018995	C0025023	638.75
C0015300	C0040165	1261.75
C0002962	C0032143	494.75
C0040038	C0039070	1226.75
C0003864	C0025587	1254
C0030232	C1883552	1389.75
C0034494	C0702166	406.25
C0232197	C0004147	1191.5
C0006840	C0392071	807.5
C0085208	C0002600	652.25
C0005367	C0039286	857.5
C0032617	C0162275	1433.25
C0553735	C0001367	603.75
C0001927	C0073992	1104
C0040034	C0018834	509.25
C0030305	C0016204	333
C0162275	C0021641	1243.5
C0019134	C0033603	1344.75
C0009262	C0032950	772.25
C0152447	C0040822	354
C0039128	C0497327	1364
C0025289	C0025287	1225.5
C0877781	C0000970	544.5
C1883552	C0017687	799
C0015772	C0051696	528
C0012963	C0030049	522
C0040038	C0232197	1148.5
C0878544	C0002962	1287.25
C0026946	C0005716	1302.75
C0006949	C0031507	797.5
C0041948	C0013911	517
C0014563	C0028351	727.25
C0035435	C0917801	379
C0242339	C0016157	1355.5
C0001911	C0025023	706.5
C0344370	C2004489	525.75
C1623038	C0002871	1187
C0039128	C0220892	1310
C0232471	C0020175	1315.75
C0003615	C0031154	1263
C0717550	C0288171	720.5
C0004153	C0858529	1179
C0019158	C0019209	1350
C0033860	C0003864	1168.75
C0235250	C0027497	1368.75
C0011175	C0013369	1299.25
C0040038	C0019134	1380.25
C0032285	C0036690	1266.25
C0085631	C0026549	1115
C0070166	C0286651	1329.75
C0007537	C0007557	1122.25
C0033860	C0054836	353.5
C0036323	C0242723	1303.75
C0553735	C0037384	305.75
C1883552	C0013911	1341.25
C0039070	C1883552	1291.5
C0232197	C0002962	1248
C0021400	C0032285	1354
C0035508	C0034642	1350.25
C0032285	C1883552	1265.75
C0028978	C0025598	652
C0220892	C0020740	358.25
C0018834	C0015620	1395.75
C0021359	C0003128	1399.5
C0010520	C0014563	710.25
C0009421	C0020456	1313.5
C0070166	C0043031	1322
C0149651	C0885057	246.25
C0002962	C0858529	1128.25
C0002871	C0060277	1375.5
C0041296	C0019079	1338.5
C0007297	C0027497	1463
C0003864	C0002726	1127.25
C0001824	C0023530	1238
C0012265	C0012373	1073.25
C0028734	C0011847	1349.75
C0011847	C0032617	1439.75
C0005747	C0270327	261
C0003864	C0035435	1340
C0011847	C0020456	1279.25
C0011603	C1998461	1258.25
C0004093	C1883552	1273
C0002600	C0016365	770
C0751229	C0037384	1252.25
C0003129	C0036572	1285
C0039070	C0002333	342.25
C0043031	C0004057	1352
C0008947	C0026196	716.25
C0020676	C0557875	1309.5
C0018021	C0020676	1424
C0022116	C0995182	318.25
C0004153	C0152447	546.25
C0019209	C0019214	1370.5
C0009214	C0027358	1209.75
C0557875	C0751229	1363.5
C0030232	C0060277	1382.75
C0002962	C0025859	1256
C0286651	C0024027	1329.75
C0065374	C0072973	753.75
C0877781	C0017887	664.5
C0014038	C0025287	1247
C0854467	C0008168	1280
C0152149	C0040460	292.25
C0007559	C0007561	1337.75
C0019112	C0021359	282.25
C0054836	C0717550	736.5
C0040485	C0037763	1377.5
C0013404	C0010520	1414.75
C0002144	C0009262	1406.5
C0030305	C0086543	345.5
C0246719	C0021641	1017.5
C0043144	C0038450	1309
C0041948	C0004057	300
C0009186	C0019655	1273
C0005740	C0012772	296.25
C0032285	C0013404	1341.5
C0020175	C0038187	1429.5
C0033687	C0011847	1439.5
C0242339	C0008402	1261.5
C0033860	C0004153	321.75
C0004096	C0451641	262.75
C0001824	C0002871	1359.5
C0003126	C0003564	1208.5
C0012833	C0042571	1398.25
C0018834	C0081876	1511
C0025289	C0018681	1483.25
C1998461	C0040485	252.25
C0040038	C0013404	1325.5
C0036494	C0149651	299.5
C0039128	C0018081	1432.5
C0007398	C0023380	1107.75
C0232197	C0002962	1368.25
C0037384	C0221232	221
C0242339	C0020473	1354.25
C0043066	C0003129	360.25
C0023570	C0006982	1575
C0878544	C0026196	358.25
C0001962	C0001975	1514.5
C0030305	C0332566	318.25
C0007557	C0007561	1295.5
C0027497	C0027498	1456.75
C0029456	C0878544	326.25
C0021359	C0003128	1452
C0033687	C0026196	319.25
C0085636	C0025287	1319.25
C0004153	C0002962	1357.75
C0028754	C0037384	1439.75
C0002940	C0029456	275.5
C0060277	C0060277	1550.5
C0019158	C0018926	1294.5
C0232955	C0232962	726.75
C0242339	C0060277	371.5
C0011847	C0162275	1394.75
C0019270	C0013456	239
C0028351	C0033487	1121
C0043031	C0995182	277.25
C0004134	C0001962	1387.25
C0011175	C0017160	1427.75
C0086543	C0027358	249
C0037763	C0016860	325.75
C0011633	C0026848	1255.25
C0038187	C0003123	1427.75
C0027497	C0061851	1479.25
C0009319	C0014544	362.75
C0206160	C0043031	329.5
C0276185	C0037384	252.5
C0235250	C0061851	1456.5
C0301532	C0039840	1347
C0242339	C0002962	1301.25
C0002871	C0060277	1469.25
C0076275	C0025598	864.5
C0018681	C0000970	1423.75
C0070166	C0060657	749
C0017160	C0013369	1409.75
C0002962	C0013404	1364
C0015300	C0020550	1470.5
C2004489	C0081876	1306
C0031154	C0004134	276.5
C0007561	C0007557	1281.75
C0018933	C0030232	752.25
C2004489	C0018834	1298.25
C0011847	C0021641	1485
C0002962	C0070166	1294.75
C0009090	C0017887	311
C0242339	C0004153	1303.25
C0022116	C0022251	1363
C0040460	C0004134	268
C1998461	C0018834	279.5
C0040038	C0043031	1353
C0025289	C0007561	1295.5
C0011847	C0085602	1459.5
C0014038	C0025289	1325.75
C0034642	C0016860	1379.5
C0015620	C0034665	1351
C0017536	C0233576	226.75
C0020676	C0040165	1473
C0232197	C0018520	293
C0006309	C0027358	297.5
C0235250	C0027498	1475.5
C0013369	C0116569	257
C0013456	C0233212	253.25
C0242339	C0286651	1425.5
C0442874	C0011847	1471.75
C0009951	C0001962	1306.25
C0030193	C0026549	1462.75
C0286651	C0074554	1436
C0024730	C0000970	241.5
C0018834	C0020740	1308.25
C0014025	C0065374	1420.5
C0043031	C0042878	1441.25
C0162275	C0038187	1363.25
C0003850	C0022116	1399.5
C0019158	C0000970	1378.75
C0920289	C0015672	1389
C0009951	C0014544	1386.75
C0497327	C0995182	215.5
C0085602	C0032617	1399.75
C0028754	C0011847	1417.25
C0032285	C0007561	1370.5
C0006644	C0039771	787.25
